// () -> l l, + -> t
// 34(1270)
module FLIPFLOP_I(
        input wire Clk,
        input wire notClk,
        input wire P2_Set_ILDrn_B,        // 0001 0000
        input wire P2_Set_ILDrn_C,        // 0001 0001
        input wire P2_Set_ILDrn_D,        // 0001 0010
        input wire P2_Set_ILDrn_E,        // 0001 0011
        input wire P2_Set_ILDrn_H,        // 0001 0100
        input wire P2_Set_ILDrn_L,        // 0001 0101
        input wire P2_Set_ILDrn_A,        // 0001 0111
        input wire P2_Set_ILDrlIXtdl_B,   // 0010 0000
        input wire P2_Set_ILDrlIXtdl_C,   // 0010 0001
        input wire P2_Set_ILDrlIXtdl_D,   // 0010 0010
        input wire P2_Set_ILDrlIXtdl_E,   // 0010 0011
        input wire P2_Set_ILDrlIXtdl_H,   // 0010 0100
        input wire P2_Set_ILDrlIXtdl_L,   // 0010 0101
        input wire P2_Set_ILDrlIXtdl_A,   // 0010 0111
        input wire P2_Set_ILDrlIYtdl_B,   // 0011 0000
        input wire P2_Set_ILDrlIYtdl_C,   // 0011 0001
        input wire P2_Set_ILDrlIYtdl_D,   // 0011 0010
        input wire P2_Set_ILDrlIYtdl_E,   // 0011 0011
        input wire P2_Set_ILDrlIYtdl_H,   // 0011 0100
        input wire P2_Set_ILDrlIYtdl_L,   // 0011 0101
        input wire P2_Set_ILDrlIYtdl_A,   // 0011 0111
        input wire P2_Set_ILDlIXtdlr_B,   // 0100 0000
        input wire P2_Set_ILDlIXtdlr_C,   // 0100 0001
        input wire P2_Set_ILDlIXtdlr_D,   // 0100 0010
        input wire P2_Set_ILDlIXtdlr_E,   // 0100 0011
        input wire P2_Set_ILDlIXtdlr_H,   // 0100 0100
        input wire P2_Set_ILDlIXtdlr_L,   // 0100 0101
        input wire P2_Set_ILDlIXtdlr_A,   // 0100 0111
        input wire P2_Set_ILDlIYtdlr_B,   // 0101 0000
        input wire P2_Set_ILDlIYtdlr_C,   // 0101 0001
        input wire P2_Set_ILDlIYtdlr_D,   // 0101 0010
        input wire P2_Set_ILDlIYtdlr_E,   // 0101 0011
        input wire P2_Set_ILDlIYtdlr_H,   // 0101 0100
        input wire P2_Set_ILDlIYtdlr_L,   // 0101 0101
        input wire P2_Set_ILDlIYtdlr_A,   // 0101 0111
        input wire P2_Set_ILDlHLln,       // 0000 0001
        input wire P2_Set_ILDlIXtdln_0,   // 1111 1010
        input wire P2_Set_ILDlIXtdln_1,   // 1111 1011
        input wire P2_Set_ILDlIYtdln_0,   // 1111 1110
        input wire P2_Set_ILDlIYtdln_1,   // 1111 1111
        input wire P2_Set_ILDAlnnl_0,     // 0000 0100
        input wire P2_Set_ILDAlnnl_1,     // 0000 0101
        input wire P2_Set_ILDlnnlA_0,     // 0000 1000
        input wire P2_Set_ILDlnnlA_1,     // 0000 1001
        input wire P2_Set_ILDddnn_BC_0,   // 0110 0000
        input wire P2_Set_ILDddnn_DE_0,   // 0110 0001
        input wire P2_Set_ILDddnn_HL_0,   // 0110 0010
        input wire P2_Set_ILDddnn_SP_0,   // 0110 0011
        input wire P2_Set_ILDddnn_BC_1,   // 0110 0100
        input wire P2_Set_ILDddnn_DE_1,   // 0110 0101
        input wire P2_Set_ILDddnn_HL_1,   // 0110 0110
        input wire P2_Set_ILDddnn_SP_1,   // 0110 0111
        input wire P2_Set_ILDIXnn_0,      // 0000 1010
        input wire P2_Set_ILDIXnn_1,      // 0000 1011
        input wire P2_Set_ILDIYnn_0,      // 0000 1110
        input wire P2_Set_ILDIYnn_1,      // 0000 1111
        input wire P2_Set_ILDHLlnnl_0,    // 0000 1100
        input wire P2_Set_ILDHLlnnl_1,    // 0000 1101
        input wire P2_Set_ILDddlnnl_BC_0, // 0111 0000
        input wire P2_Set_ILDddlnnl_DE_0, // 0111 0001
        input wire P2_Set_ILDddlnnl_HL_0, // 0111 0010
        input wire P2_Set_ILDddlnnl_SP_0, // 0111 0011
        input wire P2_Set_ILDddlnnl_BC_1, // 0111 0100
        input wire P2_Set_ILDddlnnl_DE_1, // 0111 0101
        input wire P2_Set_ILDddlnnl_HL_1, // 0111 0110
        input wire P2_Set_ILDddlnnl_SP_1, // 0111 0111
        input wire P2_Set_ILDIXlnnl_0,    // 0001 1010
        input wire P2_Set_ILDIXlnnl_1,    // 0001 1011
        input wire P2_Set_ILDIYlnnl_0,    // 0001 1110
        input wire P2_Set_ILDIYlnnl_1,    // 0001 1111
        input wire P2_Set_ILDlnnlHL_0,    // 0000 0010
        input wire P2_Set_ILDlnnlHL_1,    // 0000 0011
        input wire P2_Set_ILDlnnldd_BC_0, // 1000 0000
        input wire P2_Set_ILDlnnldd_DE_0, // 1000 0001
        input wire P2_Set_ILDlnnldd_HL_0, // 1000 0010
        input wire P2_Set_ILDlnnldd_SP_0, // 1000 0011
        input wire P2_Set_ILDlnnldd_BC_1, // 1000 0100
        input wire P2_Set_ILDlnnldd_DE_1, // 1000 0101
        input wire P2_Set_ILDlnnldd_HL_1, // 1000 0110
        input wire P2_Set_ILDlnnldd_SP_1, // 1000 0111
        input wire P2_Set_ILDlnnlIX_0,    // 0010 1010
        input wire P2_Set_ILDlnnlIX_1,    // 0010 1011
        input wire P2_Set_ILDlnnlIY_0,    // 0010 1110
        input wire P2_Set_ILDlnnlIY_1,    // 0010 1111
        input wire P2_Set_IADDAn,         // 1111 0000
        input wire P2_Set_IADDAlIXtdl,    // 1100 1000
        input wire P2_Set_IADDAlIYtdl,    // 1101 1000
        input wire P2_Set_IADCAn,         // 1111 0100
        input wire P2_Set_IADCAlIXtdl,    // 1100 1100
        input wire P2_Set_IADCAlIYtdl,    // 1101 1100
        input wire P2_Set_ISUBAn,         // 1111 0001
        input wire P2_Set_ISUBAlIXtdl,    // 1100 1001
        input wire P2_Set_ISUBAlIYtdl,    // 1101 1001
        input wire P2_Set_ISBCAn,         // 1111 0101
        input wire P2_Set_ISBCAlIXtdl,    // 1100 1101
        input wire P2_Set_ISBCAlIYtdl,    // 1101 1101
        input wire P2_Set_IANDn,          // 1111 0010
        input wire P2_Set_IANDlIXtdl,     // 1100 1010
        input wire P2_Set_IANDlIYtdl,     // 1101 1010
        input wire P2_Set_IORn,           // 1111 0011
        input wire P2_Set_IORlIXtdl,      // 1100 1011
        input wire P2_Set_IORlIYtdl,      // 1101 1011
        input wire P2_Set_IXORn,          // 1111 0110
        input wire P2_Set_IXORlIXtdl,     // 1100 1110
        input wire P2_Set_IXORlIYtdl,     // 1101 1110
        input wire P2_Set_ICPn,           // 1111 0111
        input wire P2_Set_ICPlIXtdl,      // 1100 1111
        input wire P2_Set_ICPlIYtdl,      // 1101 1111
        input wire P2_Set_IINClIXtdl,     // 1111 1000
        input wire P2_Set_IINClIYtdl,     // 1111 1001
        input wire P2_Set_IDEClIXtdl,     // 1111 1100
        input wire P2_Set_IDEClIYtdl,     // 1111 1101
        input wire P2_Set_IJPnn_0,        // 0000 0110
        input wire P2_Set_IJPnn_1,        // 0000 0111
        input wire P2_Set_IJPccnn_0_0,    // 0100 1000
        input wire P2_Set_IJPccnn_1_0,    // 0100 1001
        input wire P2_Set_IJPccnn_2_0,    // 0100 1010
        input wire P2_Set_IJPccnn_3_0,    // 0100 1011
        input wire P2_Set_IJPccnn_4_0,    // 0100 1100
        input wire P2_Set_IJPccnn_5_0,    // 0100 1101
        input wire P2_Set_IJPccnn_6_0,    // 0100 1110
        input wire P2_Set_IJPccnn_7_0,    // 0100 1111
        input wire P2_Set_IJPccnn_0_1,    // 0101 1000
        input wire P2_Set_IJPccnn_1_1,    // 0101 1001
        input wire P2_Set_IJPccnn_2_1,    // 0101 1010
        input wire P2_Set_IJPccnn_3_1,    // 0101 1011
        input wire P2_Set_IJPccnn_4_1,    // 0101 1100
        input wire P2_Set_IJPccnn_5_1,    // 0101 1101
        input wire P2_Set_IJPccnn_6_1,    // 0101 1110
        input wire P2_Set_IJPccnn_7_1,    // 0101 1111
        input wire P2_Set_IJRe,           // 0011 1000
        input wire P2_Set_IJRCe,          // 0011 1010
        input wire P2_Set_IJRNCe,         // 0011 1011
        input wire P2_Set_IJRZe,          // 0011 1110
        input wire P2_Set_IJRNZe,         // 0011 1111
        input wire P2_Set_IDJNZe,         // 0011 1100
        input wire P2_Set_ICALLnn_0,      // 0001 1100
        input wire P2_Set_ICALLnn_1,      // 0001 1101
        input wire P2_Set_IINAlnl,        // 0010 1000
        input wire P2_Set_IOUTlnlA,       // 0010 1001
        input wire P2_Set_ICALLnn_0_0,    // 1000 1000
        input wire P2_Set_ICALLnn_1_0,    // 1000 1001
        input wire P2_Set_ICALLnn_2_0,    // 1000 1010
        input wire P2_Set_ICALLnn_3_0,    // 1000 1011
        input wire P2_Set_ICALLnn_4_0,    // 1000 1100
        input wire P2_Set_ICALLnn_5_0,    // 1000 1101
        input wire P2_Set_ICALLnn_6_0,    // 1000 1110
        input wire P2_Set_ICALLnn_7_0,    // 1000 1111
        input wire P2_Set_ICALLnn_0_1,    // 1001 1000
        input wire P2_Set_ICALLnn_1_1,    // 1001 1001
        input wire P2_Set_ICALLnn_2_1,    // 1001 1010
        input wire P2_Set_ICALLnn_3_1,    // 1001 1011
        input wire P2_Set_ICALLnn_4_1,    // 1001 1100
        input wire P2_Set_ICALLnn_5_1,    // 1001 1101
        input wire P2_Set_ICALLnn_6_1,    // 1001 1110
        input wire P2_Set_ICALLnn_7_1,    // 1001 1111
        input wire P2_Reset_ITABLE,
        input wire P2_Reset_ALLUNOFFICIALFF,
        // 7654 3210
        output wire [7:0] ITABLE,
        output wire [7:0] notITABLE
    );

    // wire notClk = ~Clk;

    wire _encoded0;
    wire _encoded1;
    wire _encoded2;
    wire _encoded3;
    wire _encoded4;
    wire _encoded5;
    wire _encoded6;
    wire _encoded7;

    //
    // encode
    //

    FLIPFLOP_I_encoder_0 encoder0(
        .P2_Set_ILDrn_C(P2_Set_ILDrn_C),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIXtdl_C(P2_Set_ILDrlIXtdl_C),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdlr_C(P2_Set_ILDlIXtdlr_C),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlHLln(P2_Set_ILDlHLln),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDAlnnl_1(P2_Set_ILDAlnnl_1),
        .P2_Set_ILDlnnlA_1(P2_Set_ILDlnnlA_1),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnlHL_1(P2_Set_ILDlnnlHL_1),
        .P2_Set_ILDlnnldd_DE_0(P2_Set_ILDlnnldd_DE_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Set_ICALLnn_1_0(P2_Set_ICALLnn_1_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLnn_3_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLnn_5_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLnn_1_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .encoded0(_encoded0)
    );

    FLIPFLOP_I_encoder_1 encoder1(
        .P2_Set_ILDrn_D(P2_Set_ILDrn_D),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIXtdl_D(P2_Set_ILDrlIXtdl_D),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdlr_D(P2_Set_ILDlIXtdlr_D),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDIXnn_0(P2_Set_ILDIXnn_0),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnlHL_0(P2_Set_ILDlnnlHL_0),
        .P2_Set_ILDlnnlHL_1(P2_Set_ILDlnnlHL_1),
        .P2_Set_ILDlnnldd_HL_0(P2_Set_ILDlnnldd_HL_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IJPnn_0(P2_Set_IJPnn_0),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_ICALLnn_2_0(P2_Set_ICALLnn_2_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLnn_3_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .encoded1(_encoded1)
    );

    FLIPFLOP_I_encoder_2 encoder2(
        .P2_Set_ILDrn_H(P2_Set_ILDrn_H),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIXtdl_H(P2_Set_ILDrlIXtdl_H),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdlr_H(P2_Set_ILDlIXtdlr_H),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDAlnnl_0(P2_Set_ILDAlnnl_0),
        .P2_Set_ILDAlnnl_1(P2_Set_ILDAlnnl_1),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDHLlnnl_0(P2_Set_ILDHLlnnl_0),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnldd_BC_1(P2_Set_ILDlnnldd_BC_1),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPnn_0(P2_Set_IJPnn_0),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_ICALLnn_4_0(P2_Set_ICALLnn_4_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLnn_5_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .encoded2(_encoded2)
    );

    FLIPFLOP_I_encoder_3 encoder3(
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDlnnlA_0(P2_Set_ILDlnnlA_0),
        .P2_Set_ILDlnnlA_1(P2_Set_ILDlnnlA_1),
        .P2_Set_ILDIXnn_0(P2_Set_ILDIXnn_0),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDHLlnnl_0(P2_Set_ILDHLlnnl_0),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPccnn_0_0(P2_Set_IJPccnn_0_0),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_IINAlnl(P2_Set_IINAlnl),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Set_ICALLnn_0_0(P2_Set_ICALLnn_0_0),
        .P2_Set_ICALLnn_1_0(P2_Set_ICALLnn_1_0),
        .P2_Set_ICALLnn_2_0(P2_Set_ICALLnn_2_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLnn_3_0),
        .P2_Set_ICALLnn_4_0(P2_Set_ICALLnn_4_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLnn_5_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_0_1(P2_Set_ICALLnn_0_1),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLnn_1_1),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .encoded3(_encoded3)
    );

    FLIPFLOP_I_encoder_4 encoder4(
        .P2_Set_ILDrn_B(P2_Set_ILDrn_B),
        .P2_Set_ILDrn_C(P2_Set_ILDrn_C),
        .P2_Set_ILDrn_D(P2_Set_ILDrn_D),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_H(P2_Set_ILDrn_H),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIYtdl_B(P2_Set_ILDrlIYtdl_B),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIYtdlr_B(P2_Set_ILDlIYtdlr_B),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_ICALLnn_0_1(P2_Set_ICALLnn_0_1),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLnn_1_1),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .encoded4(_encoded4)
    );

    FLIPFLOP_I_encoder_5 encoder5(
        .P2_Set_ILDrlIXtdl_B(P2_Set_ILDrlIXtdl_B),
        .P2_Set_ILDrlIXtdl_C(P2_Set_ILDrlIXtdl_C),
        .P2_Set_ILDrlIXtdl_D(P2_Set_ILDrlIXtdl_D),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_H(P2_Set_ILDrlIXtdl_H),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_B(P2_Set_ILDrlIYtdl_B),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDddnn_BC_0(P2_Set_ILDddnn_BC_0),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IINAlnl(P2_Set_IINAlnl),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .encoded5(_encoded5)
    );

    FLIPFLOP_I_encoder_6 encoder6(
        .P2_Set_ILDlIXtdlr_B(P2_Set_ILDlIXtdlr_B),
        .P2_Set_ILDlIXtdlr_C(P2_Set_ILDlIXtdlr_C),
        .P2_Set_ILDlIXtdlr_D(P2_Set_ILDlIXtdlr_D),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_H(P2_Set_ILDlIXtdlr_H),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_B(P2_Set_ILDlIYtdlr_B),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDddnn_BC_0(P2_Set_ILDddnn_BC_0),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPccnn_0_0(P2_Set_IJPccnn_0_0),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .encoded6(_encoded6)
    );

    FLIPFLOP_I_encoder_7 encoder7(
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDlnnldd_BC_0(P2_Set_ILDlnnldd_BC_0),
        .P2_Set_ILDlnnldd_DE_0(P2_Set_ILDlnnldd_DE_0),
        .P2_Set_ILDlnnldd_HL_0(P2_Set_ILDlnnldd_HL_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDlnnldd_BC_1(P2_Set_ILDlnnldd_BC_1),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_ICALLnn_0_0(P2_Set_ICALLnn_0_0),
        .P2_Set_ICALLnn_1_0(P2_Set_ICALLnn_1_0),
        .P2_Set_ICALLnn_2_0(P2_Set_ICALLnn_2_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLnn_3_0),
        .P2_Set_ICALLnn_4_0(P2_Set_ICALLnn_4_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLnn_5_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_0_1(P2_Set_ICALLnn_0_1),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLnn_1_1),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .encoded7(_encoded7)
    );

    //
    // or
    //

    wire _not_write_0 = P2_Reset_ITABLE ~| P2_Reset_ALLUNOFFICIALFF;
    wire _not_write_1 = _encoded0 ~| _encoded1;
    wire _not_write_2 = _encoded2 ~| _encoded3;
    wire _not_write_3 = _encoded4 ~| _encoded5;
    wire _not_write_4 = _encoded6 ~| _encoded7;

    wire _write_0 = _not_write_0 ~| _not_write_0;
    wire _write_1 = _not_write_1 ~| _not_write_1;
    wire _write_2 = _not_write_2 ~| _not_write_2;
    wire _write_3 = _not_write_3 ~| _not_write_3;
    wire _write_4 = _not_write_4 ~| _not_write_4;

    wire _not_write_5 = _write_0 ~| _write_1;
    wire _write_5 = _not_write_5 ~| _not_write_5;
    wire _not_write_6 = _write_2 ~| _write_5;
    wire _write_6 = _not_write_6 ~| _not_write_6;
    wire _not_write_7 = _write_3 ~| _write_6;
    wire _write_7 = _not_write_7 ~| _not_write_7;
    wire _not_write = _write_4 ~| _write_7;
    wire _write = _not_write ~| _not_write;

    // and

    wire _ITABLE_new_ITABLE0 = notITABLE[0] ~| _write;
    wire _ITABLE_new_ITABLE1 = notITABLE[1] ~| _write;
    wire _ITABLE_new_ITABLE2 = notITABLE[2] ~| _write;
    wire _ITABLE_new_ITABLE3 = notITABLE[3] ~| _write;
    wire _ITABLE_new_ITABLE4 = notITABLE[4] ~| _write;
    wire _ITABLE_new_ITABLE5 = notITABLE[5] ~| _write;
    wire _ITABLE_new_ITABLE6 = notITABLE[6] ~| _write;
    wire _ITABLE_new_ITABLE7 = notITABLE[7] ~| _write;

    // or

    wire _ITABLE_new_not0 = _encoded0 ~| _ITABLE_new_ITABLE0;
    wire _ITABLE_new_not1 = _encoded1 ~| _ITABLE_new_ITABLE1;
    wire _ITABLE_new_not2 = _encoded2 ~| _ITABLE_new_ITABLE2;
    wire _ITABLE_new_not3 = _encoded3 ~| _ITABLE_new_ITABLE3;
    wire _ITABLE_new_not4 = _encoded4 ~| _ITABLE_new_ITABLE4;
    wire _ITABLE_new_not5 = _encoded5 ~| _ITABLE_new_ITABLE5;
    wire _ITABLE_new_not6 = _encoded6 ~| _ITABLE_new_ITABLE6;
    wire _ITABLE_new_not7 = _encoded7 ~| _ITABLE_new_ITABLE7;

    FLIPFLOP_dff itable0(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not0),
        .Q(ITABLE[0]),
        .notQ(notITABLE[0])
    );

    FLIPFLOP_dff itable1(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not1),
        .Q(ITABLE[1]),
        .notQ(notITABLE[1])
    );

    FLIPFLOP_dff itable2(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not2),
        .Q(ITABLE[2]),
        .notQ(notITABLE[2])
    );

    FLIPFLOP_dff itable3(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not3),
        .Q(ITABLE[3]),
        .notQ(notITABLE[3])
    );

    FLIPFLOP_dff itable4(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not4),
        .Q(ITABLE[4]),
        .notQ(notITABLE[4])
    );

    FLIPFLOP_dff itable5(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not5),
        .Q(ITABLE[5]),
        .notQ(notITABLE[5])
    );

    FLIPFLOP_dff itable6(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not6),
        .Q(ITABLE[6]),
        .notQ(notITABLE[6])
    );

    FLIPFLOP_dff itable7(
        .Clk(Clk),
        .notClk(notClk),
        .notD(_ITABLE_new_not7),
        .Q(ITABLE[7]),
        .notQ(notITABLE[7])
    );

endmodule