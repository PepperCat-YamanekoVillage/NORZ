// (1708)
module FLIPFLOP(
        input wire Clk,
        input wire notClk,
        input wire P2_Set_IFF1,
        input wire P2_Set_IFF2,
        input wire P2_Reset_IFF1,
        input wire P2_Reset_IFF2,
        input wire P2_EvacuateIFF,
        input wire P2_RestoreIFF,
        input wire P2_IM0,
        input wire P2_IM1,
        input wire P2_IM2,
        input wire INT,
        input wire NMI,
        input wire RESET,
        input wire WAIT,
        input wire P2_Reset_TINT,
        input wire P2_Reset_TNMI,
        input wire P2_Reset_TRSET,
        input wire P2_Set_LHALT,
        input wire P2_Reset_LHALT,
        input wire P2_Set_CM1,
        input wire P2_Set_CMR,
        input wire P2_Set_CMA,
        input wire P2_Set_CBUSRQ,
        input wire P2_Set_CRESET,
        input wire P2_Set_CNMI,
        input wire P2_Set_CINT0,
        input wire P2_Set_CINT0_RST,
        input wire P2_Set_CINT0_CALL,
        input wire P2_Set_CINT1,
        input wire P2_Set_CINT2,
        input wire P2_Reset_CM1,
        input wire P2_Reset_CMR,
        input wire P2_Reset_CMA,
        input wire P2_Reset_CBUSRQ,
        input wire P2_Reset_CRESET,
        input wire P2_Reset_CNMI,
        input wire P2_Reset_CINT,
        input wire P2_Set_XIX,
        input wire P2_Set_XIX4_0,
        input wire P2_Set_XIX4_1,
        input wire P2_Set_XIY,
        input wire P2_Set_XIY4_0,
        input wire P2_Set_XIY4_1,
        input wire P2_Set_XOTR,
        input wire P2_Set_XBIT,
        input wire P2_Reset_XIX,
        input wire P2_Reset_XIX4,
        input wire P2_Reset_XIY,
        input wire P2_Reset_XIY4,
        input wire P2_Reset_XOTR,
        input wire P2_Reset_XBIT,
        input wire P2_Set_ILDrn_B,
        input wire P2_Set_ILDrn_C,
        input wire P2_Set_ILDrn_D,
        input wire P2_Set_ILDrn_E,
        input wire P2_Set_ILDrn_H,
        input wire P2_Set_ILDrn_L,
        input wire P2_Set_ILDrn_A,
        input wire P2_Set_ILDrlIXtdl_B,
        input wire P2_Set_ILDrlIXtdl_C,
        input wire P2_Set_ILDrlIXtdl_D,
        input wire P2_Set_ILDrlIXtdl_E,
        input wire P2_Set_ILDrlIXtdl_H,
        input wire P2_Set_ILDrlIXtdl_L,
        input wire P2_Set_ILDrlIXtdl_A,
        input wire P2_Set_ILDrlIYtdl_B,
        input wire P2_Set_ILDrlIYtdl_C,
        input wire P2_Set_ILDrlIYtdl_D,
        input wire P2_Set_ILDrlIYtdl_E,
        input wire P2_Set_ILDrlIYtdl_H,
        input wire P2_Set_ILDrlIYtdl_L,
        input wire P2_Set_ILDrlIYtdl_A,
        input wire P2_Set_ILDlIXtdlr_B,
        input wire P2_Set_ILDlIXtdlr_C,
        input wire P2_Set_ILDlIXtdlr_D,
        input wire P2_Set_ILDlIXtdlr_E,
        input wire P2_Set_ILDlIXtdlr_H,
        input wire P2_Set_ILDlIXtdlr_L,
        input wire P2_Set_ILDlIXtdlr_A,
        input wire P2_Set_ILDlIYtdlr_B,
        input wire P2_Set_ILDlIYtdlr_C,
        input wire P2_Set_ILDlIYtdlr_D,
        input wire P2_Set_ILDlIYtdlr_E,
        input wire P2_Set_ILDlIYtdlr_H,
        input wire P2_Set_ILDlIYtdlr_L,
        input wire P2_Set_ILDlIYtdlr_A,
        input wire P2_Set_ILDlHLln,
        input wire P2_Set_ILDlIXtdln_0,
        input wire P2_Set_ILDlIXtdln_1,
        input wire P2_Set_ILDlIYtdln_0,
        input wire P2_Set_ILDlIYtdln_1,
        input wire P2_Set_ILDAlnnl_0,
        input wire P2_Set_ILDAlnnl_1,
        input wire P2_Set_ILDlnnlA_0,
        input wire P2_Set_ILDlnnlA_1,
        input wire P2_Set_ILDddnn_BC_0,
        input wire P2_Set_ILDddnn_DE_0,
        input wire P2_Set_ILDddnn_HL_0,
        input wire P2_Set_ILDddnn_SP_0,
        input wire P2_Set_ILDddnn_BC_1,
        input wire P2_Set_ILDddnn_DE_1,
        input wire P2_Set_ILDddnn_HL_1,
        input wire P2_Set_ILDddnn_SP_1,
        input wire P2_Set_ILDIXnn_0,
        input wire P2_Set_ILDIXnn_1,
        input wire P2_Set_ILDIYnn_0,
        input wire P2_Set_ILDIYnn_1,
        input wire P2_Set_ILDHLlnnl_0,
        input wire P2_Set_ILDHLlnnl_1,
        input wire P2_Set_ILDddlnnl_BC_0,
        input wire P2_Set_ILDddlnnl_DE_0,
        input wire P2_Set_ILDddlnnl_HL_0,
        input wire P2_Set_ILDddlnnl_SP_0,
        input wire P2_Set_ILDddlnnl_BC_1,
        input wire P2_Set_ILDddlnnl_DE_1,
        input wire P2_Set_ILDddlnnl_HL_1,
        input wire P2_Set_ILDddlnnl_SP_1,
        input wire P2_Set_ILDIXlnnl_0,
        input wire P2_Set_ILDIXlnnl_1,
        input wire P2_Set_ILDIYlnnl_0,
        input wire P2_Set_ILDIYlnnl_1,
        input wire P2_Set_ILDlnnlHL_0,
        input wire P2_Set_ILDlnnlHL_1,
        input wire P2_Set_ILDlnnldd_BC_0,
        input wire P2_Set_ILDlnnldd_DE_0,
        input wire P2_Set_ILDlnnldd_HL_0,
        input wire P2_Set_ILDlnnldd_SP_0,
        input wire P2_Set_ILDlnnldd_BC_1,
        input wire P2_Set_ILDlnnldd_DE_1,
        input wire P2_Set_ILDlnnldd_HL_1,
        input wire P2_Set_ILDlnnldd_SP_1,
        input wire P2_Set_ILDlnnlIX_0,
        input wire P2_Set_ILDlnnlIX_1,
        input wire P2_Set_ILDlnnlIY_0,
        input wire P2_Set_ILDlnnlIY_1,
        input wire P2_Set_IADDAn,
        input wire P2_Set_IADDAlIXtdl,
        input wire P2_Set_IADDAlIYtdl,
        input wire P2_Set_IADCAn,
        input wire P2_Set_IADCAlIXtdl,
        input wire P2_Set_IADCAlIYtdl,
        input wire P2_Set_ISUBAn,
        input wire P2_Set_ISUBAlIXtdl,
        input wire P2_Set_ISUBAlIYtdl,
        input wire P2_Set_ISBCAn,
        input wire P2_Set_ISBCAlIXtdl,
        input wire P2_Set_ISBCAlIYtdl,
        input wire P2_Set_IANDn,
        input wire P2_Set_IANDlIXtdl,
        input wire P2_Set_IANDlIYtdl,
        input wire P2_Set_IORn,
        input wire P2_Set_IORlIXtdl,
        input wire P2_Set_IORlIYtdl,
        input wire P2_Set_IXORn,
        input wire P2_Set_IXORlIXtdl,
        input wire P2_Set_IXORlIYtdl,
        input wire P2_Set_ICPn,
        input wire P2_Set_ICPlIXtdl,
        input wire P2_Set_ICPlIYtdl,
        input wire P2_Set_IINClIXtdl,
        input wire P2_Set_IINClIYtdl,
        input wire P2_Set_IDEClIXtdl,
        input wire P2_Set_IDEClIYtdl,
        input wire P2_Set_IJPnn_0,
        input wire P2_Set_IJPnn_1,
        input wire P2_Set_IJPccnn_0_0,
        input wire P2_Set_IJPccnn_1_0,
        input wire P2_Set_IJPccnn_2_0,
        input wire P2_Set_IJPccnn_3_0,
        input wire P2_Set_IJPccnn_4_0,
        input wire P2_Set_IJPccnn_5_0,
        input wire P2_Set_IJPccnn_6_0,
        input wire P2_Set_IJPccnn_7_0,
        input wire P2_Set_IJPccnn_0_1,
        input wire P2_Set_IJPccnn_1_1,
        input wire P2_Set_IJPccnn_2_1,
        input wire P2_Set_IJPccnn_3_1,
        input wire P2_Set_IJPccnn_4_1,
        input wire P2_Set_IJPccnn_5_1,
        input wire P2_Set_IJPccnn_6_1,
        input wire P2_Set_IJPccnn_7_1,
        input wire P2_Set_IJRe,
        input wire P2_Set_IJRCe,
        input wire P2_Set_IJRNCe,
        input wire P2_Set_IJRZe,
        input wire P2_Set_IJRNZe,
        input wire P2_Set_IDJNZe,
        input wire P2_Set_ICALLnn_0,
        input wire P2_Set_ICALLnn_1,
        input wire P2_Set_ICALLnn_0_0,
        input wire P2_Set_ICALLnn_1_0,
        input wire P2_Set_ICALLnn_2_0,
        input wire P2_Set_ICALLnn_3_0,
        input wire P2_Set_ICALLnn_4_0,
        input wire P2_Set_ICALLnn_5_0,
        input wire P2_Set_ICALLnn_6_0,
        input wire P2_Set_ICALLnn_7_0,
        input wire P2_Set_ICALLnn_0_1,
        input wire P2_Set_ICALLnn_1_1,
        input wire P2_Set_ICALLnn_2_1,
        input wire P2_Set_ICALLnn_3_1,
        input wire P2_Set_ICALLnn_4_1,
        input wire P2_Set_ICALLnn_5_1,
        input wire P2_Set_ICALLnn_6_1,
        input wire P2_Set_ICALLnn_7_1,
        input wire P2_Set_IINAlnl,
        input wire P2_Set_IOUTlnlA,
        input wire P2_Reset_ITABLE,
        input wire P2_Reset_ALLUNOFFICIALFF,
        output wire notIFF1,
        output wire IFF2,
        output wire IMFa,
        output wire IMFb,
        output wire TINT,
        output wire TNMI,
        output wire TRESET,
        output wire TWAIT,
        output wire notLHALT,
        output wire notCM1,
        output wire notCMR,
        output wire notCMA,
        output wire notCBUSRQ,
        output wire notCRESET,
        output wire notCNMI,
        output wire notCINT0,
        output wire notCINT0_RST,
        output wire notCINT0_CALL,
        output wire notCINT1,
        output wire notCINT2,
        output wire XIX,
        output wire XIX4_0,
        output wire XIX4_1,
        output wire XIY,
        output wire XIY4_0,
        output wire XIY4_1,
        output wire XOTR,
        output wire XBIT,
        output wire notXIX,
        output wire notXIX4_0,
        output wire notXIX4_1,
        output wire notXIY,
        output wire notXIY4_0,
        output wire notXIY4_1,
        output wire notXOTR,
        output wire notXBIT,
        output wire [7:0] ITABLE,
        output wire [7:0] notITABLE
    );

    FLIPFLOP_IFF iff(
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_IFF1(P2_Set_IFF1),
        .P2_Set_IFF2(P2_Set_IFF2),
        .P2_Reset_IFF1(P2_Reset_IFF1),
        .P2_Reset_IFF2(P2_Reset_IFF2),
        .P2_EvacuateIFF(P2_EvacuateIFF),
        .P2_RestoreIFF(P2_RestoreIFF),
        .notIFF1(notIFF1),
        .IFF2(IFF2)
    );

    FLIPFLOP_IMF imf(
        .Clk(Clk),
        .notClk(notClk),
        .P2_IM0(P2_IM0),
        .P2_IM1(P2_IM1),
        .P2_IM2(P2_IM2),
        .IMFa(IMFa),
        .IMFb(IMFb)
    );

    FLIPFLOP_T t(
        .Clk(Clk),
        .notClk(notClk),
        .INT(INT),
        .NMI(NMI),
        .RESET(RESET),
        .WAIT(WAIT),
        .notIFF1(notIFF1),
        .P2_Reset_TINT(P2_Reset_TINT),
        .P2_Reset_TNMI(P2_Reset_TNMI),
        .P2_Reset_TRSET(P2_Reset_TRSET),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALLUNOFFICIALFF),
        .TINT(TINT),
        .TNMI(TNMI),
        .TRESET(TRESET),
        .TWAIT(TWAIT)
    );

    FLIPFLOP_L l(
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_LHALT(P2_Set_LHALT),
        .P2_Reset_LHALT(P2_Reset_LHALT),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALLUNOFFICIALFF),
        .notLHALT(notLHALT)
    );

    FLIPFLOP_C c(
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_CM1(P2_Set_CM1),
        .P2_Set_CMR(P2_Set_CMR),
        .P2_Set_CMA(P2_Set_CMA),
        .P2_Set_CBUSRQ(P2_Set_CBUSRQ),
        .P2_Set_CRESET(P2_Set_CRESET),
        .P2_Set_CNMI(P2_Set_CNMI),
        .P2_Set_CINT0(P2_Set_CINT0),
        .P2_Set_CINT0_RST(P2_Set_CINT0_RST),
        .P2_Set_CINT0_CALL(P2_Set_CINT0_CALL),
        .P2_Set_CINT1(P2_Set_CINT1),
        .P2_Set_CINT2(P2_Set_CINT2),
        .P2_Reset_CM1(P2_Reset_CM1),
        .P2_Reset_CMR(P2_Reset_CMR),
        .P2_Reset_CMA(P2_Reset_CMA),
        .P2_Reset_CBUSRQ(P2_Reset_CBUSRQ),
        .P2_Reset_CRESET(P2_Reset_CRESET),
        .P2_Reset_CNMI(P2_Reset_CNMI),
        .P2_Reset_CINT(P2_Reset_CINT),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALLUNOFFICIALFF),
        .notCM1(notCM1),
        .notCMR(notCMR),
        .notCMA(notCMA),
        .notCBUSRQ(notCBUSRQ),
        .notCRESET(notCRESET),
        .notCNMI(notCNMI),
        .notCINT0(notCINT0),
        .notCINT0_RST(notCINT0_RST),
        .notCINT0_CALL(notCINT0_CALL),
        .notCINT1(notCINT1),
        .notCINT2(notCINT2)
    );

    FLIPFLOP_X x(
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_XIX(P2_Set_XIX),
        .P2_Set_XIX4_0(P2_Set_XIX4_0),
        .P2_Set_XIX4_1(P2_Set_XIX4_1),
        .P2_Set_XIY(P2_Set_XIY),
        .P2_Set_XIY4_0(P2_Set_XIY4_0),
        .P2_Set_XIY4_1(P2_Set_XIY4_1),
        .P2_Set_XOTR(P2_Set_XOTR),
        .P2_Set_XBIT(P2_Set_XBIT),
        .P2_Reset_XIX(P2_Reset_XIX),
        .P2_Reset_XIX4(P2_Reset_XIX4),
        .P2_Reset_XIY(P2_Reset_XIY),
        .P2_Reset_XIY4(P2_Reset_XIY4),
        .P2_Reset_XOTR(P2_Reset_XOTR),
        .P2_Reset_XBIT(P2_Reset_XBIT),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALLUNOFFICIALFF),
        .XIX(XIX),
        .XIX4_0(XIX4_0),
        .XIX4_1(XIX4_1),
        .XIY(XIY),
        .XIY4_0(XIY4_0),
        .XIY4_1(XIY4_1),
        .XOTR(XOTR),
        .XBIT(XBIT),
        .notXIX(notXIX),
        .notXIX4_0(notXIX4_0),
        .notXIX4_1(notXIX4_1),
        .notXIY(notXIY),
        .notXIY4_0(notXIY4_0),
        .notXIY4_1(notXIY4_1),
        .notXOTR(notXOTR),
        .notXBIT(notXBIT)
    );

    FLIPFLOP_I i(
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_ILDrn_B(P2_Set_ILDrn_B),
        .P2_Set_ILDrn_C(P2_Set_ILDrn_C),
        .P2_Set_ILDrn_D(P2_Set_ILDrn_D),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_H(P2_Set_ILDrn_H),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIXtdl_B(P2_Set_ILDrlIXtdl_B),
        .P2_Set_ILDrlIXtdl_C(P2_Set_ILDrlIXtdl_C),
        .P2_Set_ILDrlIXtdl_D(P2_Set_ILDrlIXtdl_D),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_H(P2_Set_ILDrlIXtdl_H),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_B(P2_Set_ILDrlIYtdl_B),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdlr_B(P2_Set_ILDlIXtdlr_B),
        .P2_Set_ILDlIXtdlr_C(P2_Set_ILDlIXtdlr_C),
        .P2_Set_ILDlIXtdlr_D(P2_Set_ILDlIXtdlr_D),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_H(P2_Set_ILDlIXtdlr_H),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_B(P2_Set_ILDlIYtdlr_B),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlHLln(P2_Set_ILDlHLln),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDAlnnl_0(P2_Set_ILDAlnnl_0),
        .P2_Set_ILDAlnnl_1(P2_Set_ILDAlnnl_1),
        .P2_Set_ILDlnnlA_0(P2_Set_ILDlnnlA_0),
        .P2_Set_ILDlnnlA_1(P2_Set_ILDlnnlA_1),
        .P2_Set_ILDddnn_BC_0(P2_Set_ILDddnn_BC_0),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDIXnn_0(P2_Set_ILDIXnn_0),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDHLlnnl_0(P2_Set_ILDHLlnnl_0),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnlHL_0(P2_Set_ILDlnnlHL_0),
        .P2_Set_ILDlnnlHL_1(P2_Set_ILDlnnlHL_1),
        .P2_Set_ILDlnnldd_BC_0(P2_Set_ILDlnnldd_BC_0),
        .P2_Set_ILDlnnldd_DE_0(P2_Set_ILDlnnldd_DE_0),
        .P2_Set_ILDlnnldd_HL_0(P2_Set_ILDlnnldd_HL_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDlnnldd_BC_1(P2_Set_ILDlnnldd_BC_1),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPnn_0(P2_Set_IJPnn_0),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .P2_Set_IJPccnn_0_0(P2_Set_IJPccnn_0_0),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_IINAlnl(P2_Set_IINAlnl),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Set_ICALLnn_0_0(P2_Set_ICALLnn_0_0),
        .P2_Set_ICALLnn_1_0(P2_Set_ICALLnn_1_0),
        .P2_Set_ICALLnn_2_0(P2_Set_ICALLnn_2_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLnn_3_0),
        .P2_Set_ICALLnn_4_0(P2_Set_ICALLnn_4_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLnn_5_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLnn_7_0),
        .P2_Set_ICALLnn_0_1(P2_Set_ICALLnn_0_1),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLnn_1_1),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLnn_3_1),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLnn_7_1),
        .P2_Reset_ITABLE(P2_Reset_ITABLE),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALLUNOFFICIALFF),
        .ITABLE(ITABLE),
        .notITABLE(notITABLE)
    );

endmodule