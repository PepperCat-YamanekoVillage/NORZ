// 107(13740)
module NORZ(
        output wire [15:0] interfaceAd,
        // 本当はinterfaceDt_inとinterfaceDt_outはinoutで同一だけどdigitalJSがエラーおこすので分けている
        input wire [7:0] interfaceDt_in,
        output wire [7:0] interfaceDt_out,
        input wire BUSRQ,
        output wire interfaceBUSAK,
        output wire interfaceMREQ,
        output wire interfaceRD,
        output wire interfaceWR,
        output wire interfaceRFSH,
        output wire interfaceIORQ,
        output wire interfaceM1,
        input wire RESET,
        input wire WAIT,
        output wire interfaceHALT,
        input wire NMI,
        input wire INT,
        input wire Clk,
        // input wire VCC,
        // input wire GND,
        //
        // for debug
        //
        output wire [7:0] _A,
        output wire [7:0] _F,
        output wire [7:0] _B,
        output wire [7:0] _C,
        output wire [7:0] _D,
        output wire [7:0] _E,
        output wire [7:0] _H,
        output wire [7:0] _L,
        output wire [15:0] _PC,
        output wire [15:0] _SP,
        output wire [15:0] _IX,
        output wire [15:0] _IY,
        output wire [7:0] _I,
        output wire [7:0] _Dt,
        output wire [7:0] _Dtex,
        output wire [7:0] _Dtcs,
        output wire [7:0] _OP,
        output wire [7:0] _OPold,
        output wire [7:0] _R,
        output wire [4:0] _XPT,
        output wire [7:0] _ITABLE,
        output wire [15:0] _ALU
    );

    // for debug
    assign _A = ~notA;
    assign _F = ~notF;
    assign _B = ~notB;
    assign _C = ~notC;
    assign _D = ~notD;
    assign _E = ~notE;
    assign _H = ~notH;
    assign _L = ~notL;
    assign _PC = ~notPC;
    assign _SP = ~notSP;
    assign _IX = ~notIX;
    assign _IY = ~notIY;
    assign _I = ~notI;
    assign _Dt = ~notDt;
    assign _Dtex = ~notDtex;
    assign _R = ~notR;
    assign _Dtcs = Dtcs;
    assign _OP = OP;
    assign _OPold = OPold;
    assign _XPT = XPT;
    assign _ITABLE = ITABLE;
    assign _ALU = ~notALU;

    wire notClk = Clk ~| Clk;

    wire [7:0] notA;
    wire [7:0] notF;
    wire [7:0] notB;
    wire [7:0] notC;
    wire [7:0] notD;
    wire [7:0] notE;
    wire [7:0] notH;
    wire [7:0] notL;
    wire [15:0] notPC;
    wire [15:0] notSP;
    wire [15:0] notIX;
    wire [15:0] notIY;
    wire [7:0] notI;
    wire [7:0] notDt;
    wire [7:0] notDtex;
    wire [7:0] Dtcs;
    wire [7:0] notDtcs;
    wire [7:0] OP;
    wire [7:0] notOP;
    wire [7:0] OPold;
    wire [7:0] notOPold;
    wire [7:0] notR;
    wire [4:0] XPT;
    wire [4:0] notXPT;
    wire [7:0] ITABLE;
    wire [7:0] notITABLE;
    wire [15:0] notALU;
    wire [7:0] Din;

    wire [7:0] notDin = ~Din; // 8

    ALU alu( // 1832 + 19
        .notA(notA),
        .notF(notF),
        .notB(notB),
        .notC(notC),
        .notD(notD),
        .notE(notE),
        .notH(notH),
        .notL(notL),
        .notDt(notDt),
        .notDtcs(notDtcs),
        .notDin(notDin),
        .notR(notR),
        .notI(notI),
        .notOP(notOP),
        .notOPold(notOPold),
        .notPC(notPC),
        .notSP(notSP),
        .notIX(notIX),
        .notIY(notIY),
        .Flag_C(~notF[0]),
        .notPA_Select_A_high(~PA_Select_A_high),
        .notPA_Select_B_high(~PA_Select_B_high),
        .PA_Select_C_high(PA_Select_C_high),
        .notPA_Select_D_high(~PA_Select_D_high),
        .PA_Select_E_high(PA_Select_E_high),
        .notPA_Select_H_high(~PA_Select_H_high),
        .PA_Select_L_high(PA_Select_L_high),
        .notPA_Select_Dt_high(PA_Select_Dt_high),
        .PA_Select_BC_high(PA_Select_BC_high),
        .PA_Select_DE_high(PA_Select_DE_high),
        .PA_Select_HL_high(PA_Select_HL_high),
        .notPA_Select_PC_high(PA_Select_PC_high),
        .notPA_Select_SP_high(PA_Select_SP_high),
        .notPA_Select_IX_high(PA_Select_IX_high),
        .notPA_Select_IY_high(PA_Select_IY_high),
        .PA_Select_0x1_high(0), // 未使用
        .notPA_Select_A_low(~PA_Select_A_low),
        .notPA_Select_F_low(~PA_Select_F_low),
        .notPA_Select_B_low(~PA_Select_B_low),
        .PA_Select_C_low(PA_Select_C_low),
        .notPA_Select_D_low(~PA_Select_D_low),
        .PA_Select_E_low(PA_Select_E_low),
        .notPA_Select_H_low(~PA_Select_H_low),
        .PA_Select_L_low(PA_Select_L_low),
        .notPA_Select_Dt_low(~PA_Select_Dt_low),
        .notPA_Select_Dtcs_low(~PA_Select_Dtcs_low),
        .notPA_Select_Din_low(~PA_Select_Din_low),
        .notPA_Select_R_low(~PA_Select_R_low),
        .notPA_Select_I_low(~PA_Select_I_low),
        .PA_Select_OP_low(PA_Select_OP_low),
        .PA_Select_BC_low(PA_Select_BC_low),
        .PA_Select_DE_low(PA_Select_DE_low),
        .PA_Select_HL_low(PA_Select_HL_low),
        .notPA_Select_PC_low(1), // 未使用
        .notPA_Select_SP_low(~PA_Select_SP_low),
        .notPA_Select_IX_low(~PA_Select_IX_low),
        .notPA_Select_IY_low(~PA_Select_IY_low),
        .PA_Select_IOP_low(PA_Select_IOP_low),
        .notPA_Select_OPOPold_low(~PA_Select_OPOPold_low),
        .PA_Select_0xffOP_low(PA_Select_0xffOP_low),
        .PA_Select_OPold_low(PA_Select_OPold_low),
        .PA_Select_OP_high(PA_Select_OP_high),
        .PA_Select_0x1_low(PA_Select_0x1_low),
        .PA_Select_0x8_low(PA_Select_0x8_low),
        .PA_Select_0x10_low(PA_Select_0x10_low),
        .PA_Select_0x18_low(PA_Select_0x18_low),
        .PA_Select_0x20_low(PA_Select_0x20_low),
        .PA_Select_0x28_low(PA_Select_0x28_low),
        .PA_Select_0x30_low(PA_Select_0x30_low),
        .PA_Select_0x38_low(PA_Select_0x38_low),
        .PA_Select_0x66_low(PA_Select_0x66_low),
        .PA_Select_0x99_low(PA_Select_0x99_low),
        .PA_Select_0x06_low(PA_Select_0x06_low),
        .PA_Select_0x60_low(PA_Select_0x60_low),
        .PA_Select_0x2_low(PA_Select_0x2_low),
        .PA_Select_0x4_low(PA_Select_0x4_low),
        .PA_Select_0x40_low(PA_Select_0x40_low),
        .PA_Select_0x80_low(PA_Select_0x80_low),
        .PA_NOP(PA_NOP),
        .PA_ADD(PA_ADD),
        .PA_ADC(PA_ADC),
        .PA_SUB(PA_SUB),
        .PA_SBC(PA_SBC),
        .PA_NOT(PA_NOT),
        .PA_AND(PA_AND),
        .PA_NLAND(PA_NLAND),
        .PA_OR(PA_OR),
        .PA_XOR(PA_XOR),
        .PA_RLC(PA_RLC),
        .PA_RL(PA_RL),
        .PA_SLA(PA_SLA),
        .PA_RRC(PA_RRC),
        .PA_RR(PA_RR),
        .PA_SRA(PA_SRA),
        .PA_SRL(PA_SRL),
        .PA_RLD(PA_RLD),
        .PA_RRD(PA_RRD),
        .notResult(notALU),
        .notLow0(notALULow0),
        .notLow7(notALULow7),
        .notCY4(notCY4),
        .notCY8(notCY8),
        .CY12(CY12),
        .CY16(CY16),
        .notIs8bitEqual(notIs8bitEqual),
        .is16bitEqual(is16bitEqual),
        .notIsResultLow0(notIsResultLow0),
        .isResult0(isResult0),
        .is8bitOverflow(is8bitOverflow),
        .is16bitOverflow(is16bitOverflow),
        .notIs8bitEvenParity(notIs8bitEvenParity),
        .DAA_Flag_H(DAA_Flag_H)
    );

    DECODER dec( // 5307 + 6
        .Clk(Clk),
        .notClk(notClk),
        .RESET(RESET),
        .TRESET(TRESET),
        .BUSRQ(BUSRQ),
        .TNMI(TNMI),
        .TINT(TINT),
        .notIFF1(notIFF1),
        .IMFa(IMFa),
        .IMFb(IMFb),
        .notCRESET(notCRESET),
        .notCBUSRQ(notCBUSRQ),
        .notCNMI(notCNMI),
        .notCINT0_RST(notCINT0_RST),
        .notCINT0_CALL(notCINT0_CALL),
        .notCINT0(notCINT0),
        .notCINT1(notCINT1),
        .notCINT2(notCINT2),
        .notCM1(notCM1), // XPT 0,1のみXOR
        .notCMR(notCMR), // XPT 0,1のみXOR
        .notCMA(notCMA), // XPT 0,1のみXOR
        .TWAIT(TWAIT),
        .XPT(XPT),
        .notXPT(notXPT),
        .ITABLE(ITABLE),
        .notITABLE(notITABLE),
        .OP(OP),
        .Dtcs(Dtcs),
        .notIsResultLow0(notIsResultLow0),
        .notXIX(notXIX),
        .notXIX4_0(notXIX4_0),
        .notXIX4_1(notXIX4_1),
        .notXIY(notXIY),
        .notXIY4_0(notXIY4_0),
        .notXIY4_1(notXIY4_1),
        .notXOTR(notXOTR),
        .notXBIT(notXBIT),
        .Flag_H(~notF[4]),
        .Flag_Z(~notF[6]),
        .Flag_C(~notF[0]),
        .Flag_S(~notF[7]),
        .Flag_N(~notF[1]),
        .Flag_PV(~notF[2]),
        .notFlag_Z(notF[6]),
        .P2_Set_CRESET(P2_Set_CRESET),
        .P2_Reset_ALL_except_CRESET(P2_Reset_ALL_except_CRESET),
        .P2_Set_CBUSRQ(P2_Set_CBUSRQ),
        .PI_Nullify_MREQ(PI_Nullify_MREQ),
        .PI_Nullify_RD(PI_Nullify_RD),
        .PI_Nullify_WR(PI_Nullify_WR),
        .PI_Nullify_IORQ(PI_Nullify_IORQ),
        .PI_Flag_BUSAK(PI_Flag_BUSAK),
        .PR_Halt_XPT(PR_Halt_XPT),
        .P2_Set_CNMI(P2_Set_CNMI),
        .P2_Reset_TNMI(P2_Reset_TNMI),
        .P2_Reset_LHALT(P2_Reset_LHALT),
        .P2_EvacuateIFF(P2_EvacuateIFF),
        .P2_Reset_IFF1(P2_Reset_IFF1),
        .P2_Set_CINT0(P2_Set_CINT0),
        .P2_Set_CINT1(P2_Set_CINT1),
        .P2_Set_CINT2(P2_Set_CINT2),
        .P2_Reset_TINT(P2_Reset_TINT),
        .P2_Reset_IFF2(P2_Reset_IFF2),
        .PI_Activate_Ad_high(PI_Activate_Ad_high),
        .PI_Activate_Ad_low(PI_Activate_Ad_low),
        .PI_SelectAd_PC(PI_SelectAd_PC),
        .PI_Flag_M1(PI_Flag_M1),
        .PR_Reset_XPT(PR_Reset_XPT),
        .PA_NOP(PA_NOP),
        .PR_Write_PC_low(PR_Write_PC_low),
        .PR_Write_PC_high(PR_Write_PC_high),
        .PR_Write_I(PR_Write_I),
        .PR_Write_R(PR_Write_R),
        .P2_Reset_CRESET(P2_Reset_CRESET),
        .P2_Set_CM1(P2_Set_CM1),
        .P2_IM0(P2_IM0),
        .P2_Reset_CBUSRQ(P2_Reset_CBUSRQ),
        .PR_Dec_SP(PR_Dec_SP),
        .PI_SelectDt_PC_high(PI_SelectDt_PC_high),
        .PI_SelectDt_PC_low(PI_SelectDt_PC_low),
        .PI_SelectAd_SP(PI_SelectAd_SP),
        .P2_Reset_CNMI(P2_Reset_CNMI),
        .PA_Select_0x66_low(PA_Select_0x66_low),
        .PA_Select_0x8_low(PA_Select_0x8_low),
        .PA_Select_0x10_low(PA_Select_0x10_low),
        .PA_Select_0x18_low(PA_Select_0x18_low),
        .PA_Select_0x20_low(PA_Select_0x20_low),
        .PA_Select_0x28_low(PA_Select_0x28_low),
        .PA_Select_0x30_low(PA_Select_0x30_low),
        .PA_Select_0x38_low(PA_Select_0x38_low),
        .P2_Reset_CINT(P2_Reset_CINT),
        .PA_Select_OPOPold_low(PA_Select_OPOPold_low),
        .P2_Set_CINT0_RST(P2_Set_CINT0_RST),
        .P2_Set_CINT0_CALL(P2_Set_CINT0_CALL),
        .PA_Select_IOP_low(PA_Select_IOP_low),
        .PI_Flag_IORQ(PI_Flag_IORQ),
        .PA_Select_Din_low(PA_Select_Din_low),
        .PR_Write_OP(PR_Write_OP),
        .PI_SelectAd_IR(PI_SelectAd_IR),
        .PI_Flag_RFSH(PI_Flag_RFSH),
        .PR_Inc_R(PR_Inc_R),
        .PI_Flag_MREQ(PI_Flag_MREQ),
        .PI_Flag_RD(PI_Flag_RD),
        .P2_Reset_CM1(P2_Reset_CM1),
        .PR_SlideOP(PR_SlideOP),
        .P2_Reset_CMR(P2_Reset_CMR),
        .PR_Inc_PC(PR_Inc_PC),
        .PI_Read_Dtcs(PI_Read_Dtcs),
        .PA_Select_Dtcs_low(PA_Select_Dtcs_low),
        .P2_Reset_CMA(P2_Reset_CMA),
        .PI_Flag_WR(PI_Flag_WR),
        .PI_Activate_Dt(PI_Activate_Dt),
        .PI_SelectAd_HL(PI_SelectAd_HL),
        .PI_SelectDt_OP(PI_SelectDt_OP),
        .P2_Reset_ITABLE(P2_Reset_ITABLE),
        .P2_Set_CMR(P2_Set_CMR),
        .P2_Set_ILDlnnlHL_1(P2_Set_ILDlnnlHL_1),
        .PI_SelectDt_L(PI_SelectDt_L),
        .PI_SelectDt_H(PI_SelectDt_H),
        .PI_SelectAdt1(PI_SelectAdt1),
        .PI_SelectAd_OPOPold(PI_SelectAd_OPOPold),
        .P2_Set_ILDAlnnl_1(P2_Set_ILDAlnnl_1),
        .PR_Write_A(PR_Write_A),
        .PR_InvertIn(PR_InvertIn),
        .P2_Set_CMA(P2_Set_CMA),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .PA_Select_OP_high(PA_Select_OP_high),
        .PR_Write_B(PR_Write_B),
        .PR_Write_C(PR_Write_C),
        .PR_Write_D(PR_Write_D),
        .PR_Write_E(PR_Write_E),
        .PR_Write_H(PR_Write_H),
        .PR_Write_L(PR_Write_L),
        .PA_Select_IX_high(PA_Select_IX_high),
        .PA_Select_IY_high(PA_Select_IY_high),
        .PA_Select_OP_low(PA_Select_OP_low),
        .PA_ADD(PA_ADD),
        .PR_Write_Dt(PR_Write_Dt),
        .PR_Write_Dtex(PR_Write_Dtex),
        .PI_SelectAd_DtexDt(PI_SelectAd_DtexDt),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .PR_Write_SP_low(PR_Write_SP_low),
        .PR_Write_SP_high(PR_Write_SP_high),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .PI_SelectDt_A(PI_SelectDt_A),
        .PI_SelectDt_B(PI_SelectDt_B),
        .PI_SelectDt_D(PI_SelectDt_D),
        .P2_Set_ILDlnnldd_BC_1(P2_Set_ILDlnnldd_BC_1),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .PI_SelectDt_SP_low(PI_SelectDt_SP_low),
        .PI_SelectDt_SP_high(PI_SelectDt_SP_high),
        .PA_Select_A_high(PA_Select_A_high),
        .PF_Write_S(PF_Write_S),
        .PF_Select_S_bit7(PF_Select_S_bit7),
        .PF_Write_Z(PF_Write_Z),
        .PF_Select_Z_bit24(PF_Select_Z_bit24),
        .PF_Write_H(PF_Write_H),
        .PF_Write_PV(PF_Write_PV),
        .PF_Write_N(PF_Write_N),
        .PF_Write_C(PF_Write_C),
        .PA_ADC(PA_ADC),
        .PA_SUB(PA_SUB),
        .PA_SBC(PA_SBC),
        .PA_AND(PA_AND),
        .PA_OR(PA_OR),
        .PA_XOR(PA_XOR),
        .PF_Select_H_bit22(PF_Select_H_bit22),
        .PF_Select_N_bit17(PF_Select_N_bit17),
        .PF_Select_C_bit26(PF_Select_C_bit26),
        .PF_Select_H_bit21(PF_Select_H_bit21),
        .PF_Select_C_bit23(PF_Select_C_bit23),
        .PF_Select_H_bit16(PF_Select_H_bit16), // PF_Writeで0にできる
        .PF_Select_PV_bit27(PF_Select_PV_bit27),
        .PF_Select_C_bit16(PF_Select_C_bit16), // PF_Writeで0にできる
        .PF_Select_H_bit17(PF_Select_H_bit17),
        .PF_Select_N_bit16(PF_Select_N_bit16), // PF_Writeで0にできる
        .PF_Select_PV_bit25(PF_Select_PV_bit25),
        .PR_Write_IX_low(PR_Write_IX_low),
        .PR_Write_IY_low(PR_Write_IY_low),
        .P2_Set_ILDlnnlA_1(P2_Set_ILDlnnlA_1),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .PR_Write_IX_high(PR_Write_IX_high),
        .PR_Write_IY_high(PR_Write_IY_high),
        .PI_SelectAd_AOP(PI_SelectAd_AOP),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .PI_SelectDt_IX_low(PI_SelectDt_IX_low),
        .PI_SelectDt_IY_low(PI_SelectDt_IY_low),
        .PI_SelectDt_IX_high(PI_SelectDt_IX_high),
        .PI_SelectDt_IY_high(PI_SelectDt_IY_high),
        .PA_Select_PC_high(PA_Select_PC_high),
        .PA_Select_0xffOP_low(PA_Select_0xffOP_low),
        .PA_Select_B_high(PA_Select_B_high),
        .PA_Select_0x1_low(PA_Select_0x1_low),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_ICALLccnn_0_1(P2_Set_ICALLccnn_0_1),
        .P2_Set_ICALLccnn_1_1(P2_Set_ICALLccnn_1_1),
        .P2_Set_ICALLccnn_2_1(P2_Set_ICALLccnn_2_1),
        .P2_Set_ICALLccnn_3_1(P2_Set_ICALLccnn_3_1),
        .P2_Set_ICALLccnn_4_1(P2_Set_ICALLccnn_4_1),
        .P2_Set_ICALLccnn_5_1(P2_Set_ICALLccnn_5_1),
        .P2_Set_ICALLccnn_6_1(P2_Set_ICALLccnn_6_1),
        .P2_Set_ICALLccnn_7_1(P2_Set_ICALLccnn_7_1),
        .PA_Select_Dt_high(PA_Select_Dt_high),
        .PI_SelectAd_ALU(PI_SelectAd_ALU),
        .PI_SelectDt_Dt(PI_SelectDt_Dt),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .PA_Select_OPold_low(PA_Select_OPold_low),
        .P2_Reset_XBIT(P2_Reset_XBIT),
        .PA_Select_B_low(PA_Select_B_low),
        .PA_Select_C_low(PA_Select_C_low),
        .PA_Select_D_low(PA_Select_D_low),
        .PA_Select_E_low(PA_Select_E_low),
        .PA_Select_H_low(PA_Select_H_low),
        .PA_Select_L_low(PA_Select_L_low),
        .PA_Select_A_low(PA_Select_A_low),
        .PA_Select_C_high(PA_Select_C_high),
        .PA_Select_D_high(PA_Select_D_high),
        .PA_Select_E_high(PA_Select_E_high),
        .PA_Select_H_high(PA_Select_H_high),
        .PA_Select_L_high(PA_Select_L_high),
        .PA_Select_Dt_low(PA_Select_Dt_low),
        .P2_Reset_XIX4(P2_Reset_XIX4),
        .P2_Reset_XIY4(P2_Reset_XIY4),
        .PF_Select_C_bit38(PF_Select_C_bit38),
        .PF_Select_C_bit37(PF_Select_C_bit37),
        .PA_RLC(PA_RLC),
        .PA_RL(PA_RL),
        .PA_SLA(PA_SLA),
        .PA_RRC(PA_RRC),
        .PA_RR(PA_RR),
        .PA_SRA(PA_SRA),
        .PA_SRL(PA_SRL),
        .PA_NLAND(PA_NLAND),
        .PF_Select_Z_bit40(PF_Select_Z_bit40),
        .PF_Select_Z_bit41(PF_Select_Z_bit41),
        .PF_Select_Z_bit42(PF_Select_Z_bit42),
        .PF_Select_Z_bit43(PF_Select_Z_bit43),
        .PF_Select_Z_bit44(PF_Select_Z_bit44),
        .PF_Select_Z_bit45(PF_Select_Z_bit45),
        .PF_Select_Z_bit46(PF_Select_Z_bit46),
        .PF_Select_Z_bit47(PF_Select_Z_bit47),
        .PA_Select_0x2_low(PA_Select_0x2_low),
        .PA_Select_0x4_low(PA_Select_0x4_low),
        .PA_Select_0x20_low(PA_Select_0x20_low),
        .PA_Select_0x40_low(PA_Select_0x40_low),
        .PA_Select_0x80_low(PA_Select_0x80_low),
        .P2_Set_XIX4_1(P2_Set_XIX4_1),
        .P2_Set_XIY4_1(P2_Set_XIY4_1),
        .PI_SelectAd_BC(PI_SelectAd_BC),
        .PI_SelectDt_C(PI_SelectDt_C),
        .PI_SelectDt_E(PI_SelectDt_E),
        .P2_Reset_XOTR(P2_Reset_XOTR),
        .PA_Select_HL_high(PA_Select_HL_high),
        .PF_Select_Z_bit34(PF_Select_Z_bit34),
        .PF_Select_PV_bit33(PF_Select_PV_bit33),
        .PF_Select_S_bit15(PF_Select_S_bit15),
        .PF_Select_C_bit36(PF_Select_C_bit36),
        .PF_Select_H_bit35(PF_Select_H_bit35),
        .PF_Select_C_bit32(PF_Select_C_bit32),
        .PF_Select_H_bit31(PF_Select_H_bit31),
        .PA_Select_BC_low(PA_Select_BC_low),
        .PA_Select_DE_low(PA_Select_DE_low),
        .PA_Select_HL_low(PA_Select_HL_low),
        .PA_Select_SP_low(PA_Select_SP_low),
        .P2_Set_ILDlnnldd_BC_0(P2_Set_ILDlnnldd_BC_0),
        .P2_Set_ILDlnnldd_DE_0(P2_Set_ILDlnnldd_DE_0),
        .P2_Set_ILDlnnldd_HL_0(P2_Set_ILDlnnldd_HL_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .PR_Inc_SP(PR_Inc_SP),
        .P2_RestoreIFF(P2_RestoreIFF),
        .P2_IM1(P2_IM1),
        .P2_IM2(P2_IM2),
        .PF_Select_Z_bit19(PF_Select_Z_bit19),
        .PF_Select_PV_bit18(PF_Select_PV_bit18),
        .PA_Select_I_low(PA_Select_I_low),
        .PA_Select_R_low(PA_Select_R_low),
        .PA_RRD(PA_RRD),
        .PA_RLD(PA_RLD),
        .PA_Select_BC_high(PA_Select_BC_high),
        .PF_Select_PV_bit20(PF_Select_PV_bit20),
        .PI_SelectAd_DE(PI_SelectAd_DE),
        .PA_Select_DE_high(PA_Select_DE_high),
        .P2_Reset_XIX(P2_Reset_XIX),
        .P2_Reset_XIY(P2_Reset_XIY),
        .PA_Select_IX_low(PA_Select_IX_low),
        .PA_Select_IY_low(PA_Select_IY_low),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIXnn_0(P2_Set_ILDIXnn_0),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDrlIXtdl_B(P2_Set_ILDrlIXtdl_B),
        .P2_Set_ILDrlIXtdl_C(P2_Set_ILDrlIXtdl_C),
        .P2_Set_ILDrlIXtdl_D(P2_Set_ILDrlIXtdl_D),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_H(P2_Set_ILDrlIXtdl_H),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDlIXtdlr_B(P2_Set_ILDlIXtdlr_B),
        .P2_Set_ILDlIXtdlr_C(P2_Set_ILDlIXtdlr_C),
        .P2_Set_ILDlIXtdlr_D(P2_Set_ILDlIXtdlr_D),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_H(P2_Set_ILDlIXtdlr_H),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDrlIYtdl_B(P2_Set_ILDrlIYtdl_B),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIYtdlr_B(P2_Set_ILDlIYtdlr_B),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_XIX4_0(P2_Set_XIX4_0),
        .P2_Set_XIY4_0(P2_Set_XIY4_0),
        .PI_SelectDt_Dtex(PI_SelectDt_Dtex),
        .P2_Set_LHALT(P2_Set_LHALT),
        .PR_Ex_AF_AF(PR_Ex_AF_AF),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_ILDddnn_BC_0(P2_Set_ILDddnn_BC_0),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDlnnlHL_0(P2_Set_ILDlnnlHL_0),
        .P2_Set_ILDHLlnnl_0(P2_Set_ILDHLlnnl_0),
        .P2_Set_ILDlnnlA_0(P2_Set_ILDlnnlA_0),
        .P2_Set_ILDAlnnl_0(P2_Set_ILDAlnnl_0),
        .PA_Select_SP_high(PA_Select_SP_high),
        .P2_Set_ILDrn_B(P2_Set_ILDrn_B),
        .P2_Set_ILDrn_C(P2_Set_ILDrn_C),
        .P2_Set_ILDrn_D(P2_Set_ILDrn_D),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_H(P2_Set_ILDrn_H),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDlHLln(P2_Set_ILDlHLln),
        .PA_Select_0x99_low(PA_Select_0x99_low),
        .PF_Select_S_bit23(PF_Select_S_bit23),
        .PF_Select_Z_bit21(PF_Select_Z_bit21),
        .PF_Select_C_bit29(PF_Select_C_bit29),
        .PF_Select_H_bit28(PF_Select_H_bit28),
        .PA_Select_0x60_low(PA_Select_0x60_low),
        .PA_Select_0x06_low(PA_Select_0x06_low),
        .PA_NOT(PA_NOT),
        .PF_Select_H_bit30(PF_Select_H_bit30),
        .PF_Select_C_bit0(PF_Select_C_bit0),
        .PF_Select_C_bit17(PF_Select_C_bit17),
        .PA_Select_F_low(PA_Select_F_low),
        .PR_Exx(PR_Exx),
        .PR_Write_F(PR_Write_F),
        .P2_Set_XBIT(P2_Set_XBIT),
        .PR_Ex_DE_HL(PR_Ex_DE_HL),
        .P2_Set_IFF1(P2_Set_IFF1), // <
        .P2_Set_IFF2(P2_Set_IFF2), // >
        .P2_Set_IJPccnn_0_0(P2_Set_IJPccnn_0_0),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPnn_0(P2_Set_IJPnn_0),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Set_IINAlnl(P2_Set_IINAlnl),
        .PI_SelectDt_F(PI_SelectDt_F),
        .P2_Set_ICALLccnn_0_0(P2_Set_ICALLccnn_0_0),
        .P2_Set_ICALLccnn_1_0(P2_Set_ICALLccnn_1_0),
        .P2_Set_ICALLccnn_2_0(P2_Set_ICALLccnn_2_0),
        .P2_Set_ICALLccnn_3_0(P2_Set_ICALLccnn_3_0),
        .P2_Set_ICALLccnn_4_0(P2_Set_ICALLccnn_4_0),
        .P2_Set_ICALLccnn_5_0(P2_Set_ICALLccnn_5_0),
        .P2_Set_ICALLccnn_6_0(P2_Set_ICALLccnn_6_0),
        .P2_Set_ICALLccnn_7_0(P2_Set_ICALLccnn_7_0),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_XIX(P2_Set_XIX),
        .P2_Set_XOTR(P2_Set_XOTR),
        .P2_Set_XIY(P2_Set_XIY),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_ICPn(P2_Set_ICPn)
    );

    FLIPFLOP ff( // 1708
        .Clk(Clk),
        .notClk(notClk),
        .P2_Set_IFF1(P2_Set_IFF1),
        .P2_Set_IFF2(P2_Set_IFF2),
        .P2_Reset_IFF1(P2_Reset_IFF1),
        .P2_Reset_IFF2(P2_Reset_IFF2),
        .P2_EvacuateIFF(P2_EvacuateIFF),
        .P2_RestoreIFF(P2_RestoreIFF),
        .P2_IM0(P2_IM0),
        .P2_IM1(P2_IM1),
        .P2_IM2(P2_IM2),
        .INT(INT),
        .NMI(NMI),
        .RESET(RESET),
        .WAIT(WAIT),
        .P2_Reset_TINT(P2_Reset_TINT),
        .P2_Reset_TNMI(P2_Reset_TNMI),
        .P2_Reset_TRSET(P2_Reset_TRSET),
        .P2_Set_LHALT(P2_Set_LHALT),
        .P2_Reset_LHALT(P2_Reset_LHALT),
        .P2_Set_CM1(P2_Set_CM1),
        .P2_Set_CMR(P2_Set_CMR),
        .P2_Set_CMA(P2_Set_CMA),
        .P2_Set_CBUSRQ(P2_Set_CBUSRQ),
        .P2_Set_CRESET(P2_Set_CRESET),
        .P2_Set_CNMI(P2_Set_CNMI),
        .P2_Set_CINT0(P2_Set_CINT0),
        .P2_Set_CINT0_RST(P2_Set_CINT0_RST),
        .P2_Set_CINT0_CALL(P2_Set_CINT0_CALL),
        .P2_Set_CINT1(P2_Set_CINT1),
        .P2_Set_CINT2(P2_Set_CINT2),
        .P2_Reset_CM1(P2_Reset_CM1),
        .P2_Reset_CMR(P2_Reset_CMR),
        .P2_Reset_CMA(P2_Reset_CMA),
        .P2_Reset_CBUSRQ(P2_Reset_CBUSRQ),
        .P2_Reset_CRESET(P2_Reset_CRESET),
        .P2_Reset_CNMI(P2_Reset_CNMI),
        .P2_Reset_CINT(P2_Reset_CINT),
        .P2_Set_XIX(P2_Set_XIX),
        .P2_Set_XIX4_0(P2_Set_XIX4_0),
        .P2_Set_XIX4_1(P2_Set_XIX4_1),
        .P2_Set_XIY(P2_Set_XIY),
        .P2_Set_XIY4_0(P2_Set_XIY4_0),
        .P2_Set_XIY4_1(P2_Set_XIY4_1),
        .P2_Set_XOTR(P2_Set_XOTR),
        .P2_Set_XBIT(P2_Set_XBIT),
        .P2_Reset_XIX(P2_Reset_XIX),
        .P2_Reset_XIX4(P2_Reset_XIX4),
        .P2_Reset_XIY(P2_Reset_XIY),
        .P2_Reset_XIY4(P2_Reset_XIY4),
        .P2_Reset_XOTR(P2_Reset_XOTR),
        .P2_Reset_XBIT(P2_Reset_XBIT),
        .P2_Set_ILDrn_B(P2_Set_ILDrn_B),
        .P2_Set_ILDrn_C(P2_Set_ILDrn_C),
        .P2_Set_ILDrn_D(P2_Set_ILDrn_D),
        .P2_Set_ILDrn_E(P2_Set_ILDrn_E),
        .P2_Set_ILDrn_H(P2_Set_ILDrn_H),
        .P2_Set_ILDrn_L(P2_Set_ILDrn_L),
        .P2_Set_ILDrn_A(P2_Set_ILDrn_A),
        .P2_Set_ILDrlIXtdl_B(P2_Set_ILDrlIXtdl_B),
        .P2_Set_ILDrlIXtdl_C(P2_Set_ILDrlIXtdl_C),
        .P2_Set_ILDrlIXtdl_D(P2_Set_ILDrlIXtdl_D),
        .P2_Set_ILDrlIXtdl_E(P2_Set_ILDrlIXtdl_E),
        .P2_Set_ILDrlIXtdl_H(P2_Set_ILDrlIXtdl_H),
        .P2_Set_ILDrlIXtdl_L(P2_Set_ILDrlIXtdl_L),
        .P2_Set_ILDrlIXtdl_A(P2_Set_ILDrlIXtdl_A),
        .P2_Set_ILDrlIYtdl_B(P2_Set_ILDrlIYtdl_B),
        .P2_Set_ILDrlIYtdl_C(P2_Set_ILDrlIYtdl_C),
        .P2_Set_ILDrlIYtdl_D(P2_Set_ILDrlIYtdl_D),
        .P2_Set_ILDrlIYtdl_E(P2_Set_ILDrlIYtdl_E),
        .P2_Set_ILDrlIYtdl_H(P2_Set_ILDrlIYtdl_H),
        .P2_Set_ILDrlIYtdl_L(P2_Set_ILDrlIYtdl_L),
        .P2_Set_ILDrlIYtdl_A(P2_Set_ILDrlIYtdl_A),
        .P2_Set_ILDlIXtdlr_B(P2_Set_ILDlIXtdlr_B),
        .P2_Set_ILDlIXtdlr_C(P2_Set_ILDlIXtdlr_C),
        .P2_Set_ILDlIXtdlr_D(P2_Set_ILDlIXtdlr_D),
        .P2_Set_ILDlIXtdlr_E(P2_Set_ILDlIXtdlr_E),
        .P2_Set_ILDlIXtdlr_H(P2_Set_ILDlIXtdlr_H),
        .P2_Set_ILDlIXtdlr_L(P2_Set_ILDlIXtdlr_L),
        .P2_Set_ILDlIXtdlr_A(P2_Set_ILDlIXtdlr_A),
        .P2_Set_ILDlIYtdlr_B(P2_Set_ILDlIYtdlr_B),
        .P2_Set_ILDlIYtdlr_C(P2_Set_ILDlIYtdlr_C),
        .P2_Set_ILDlIYtdlr_D(P2_Set_ILDlIYtdlr_D),
        .P2_Set_ILDlIYtdlr_E(P2_Set_ILDlIYtdlr_E),
        .P2_Set_ILDlIYtdlr_H(P2_Set_ILDlIYtdlr_H),
        .P2_Set_ILDlIYtdlr_L(P2_Set_ILDlIYtdlr_L),
        .P2_Set_ILDlIYtdlr_A(P2_Set_ILDlIYtdlr_A),
        .P2_Set_ILDlHLln(P2_Set_ILDlHLln),
        .P2_Set_ILDlIXtdln_0(P2_Set_ILDlIXtdln_0),
        .P2_Set_ILDlIXtdln_1(P2_Set_ILDlIXtdln_1),
        .P2_Set_ILDlIYtdln_0(P2_Set_ILDlIYtdln_0),
        .P2_Set_ILDlIYtdln_1(P2_Set_ILDlIYtdln_1),
        .P2_Set_ILDAlnnl_0(P2_Set_ILDAlnnl_0),
        .P2_Set_ILDAlnnl_1(P2_Set_ILDAlnnl_1),
        .P2_Set_ILDlnnlA_0(P2_Set_ILDlnnlA_0),
        .P2_Set_ILDlnnlA_1(P2_Set_ILDlnnlA_1),
        .P2_Set_ILDddnn_BC_0(P2_Set_ILDddnn_BC_0),
        .P2_Set_ILDddnn_DE_0(P2_Set_ILDddnn_DE_0),
        .P2_Set_ILDddnn_HL_0(P2_Set_ILDddnn_HL_0),
        .P2_Set_ILDddnn_SP_0(P2_Set_ILDddnn_SP_0),
        .P2_Set_ILDddnn_BC_1(P2_Set_ILDddnn_BC_1),
        .P2_Set_ILDddnn_DE_1(P2_Set_ILDddnn_DE_1),
        .P2_Set_ILDddnn_HL_1(P2_Set_ILDddnn_HL_1),
        .P2_Set_ILDddnn_SP_1(P2_Set_ILDddnn_SP_1),
        .P2_Set_ILDIXnn_0(P2_Set_ILDIXnn_0),
        .P2_Set_ILDIXnn_1(P2_Set_ILDIXnn_1),
        .P2_Set_ILDIYnn_0(P2_Set_ILDIYnn_0),
        .P2_Set_ILDIYnn_1(P2_Set_ILDIYnn_1),
        .P2_Set_ILDHLlnnl_0(P2_Set_ILDHLlnnl_0),
        .P2_Set_ILDHLlnnl_1(P2_Set_ILDHLlnnl_1),
        .P2_Set_ILDddlnnl_BC_0(P2_Set_ILDddlnnl_BC_0),
        .P2_Set_ILDddlnnl_DE_0(P2_Set_ILDddlnnl_DE_0),
        .P2_Set_ILDddlnnl_HL_0(P2_Set_ILDddlnnl_HL_0),
        .P2_Set_ILDddlnnl_SP_0(P2_Set_ILDddlnnl_SP_0),
        .P2_Set_ILDddlnnl_BC_1(P2_Set_ILDddlnnl_BC_1),
        .P2_Set_ILDddlnnl_DE_1(P2_Set_ILDddlnnl_DE_1),
        .P2_Set_ILDddlnnl_HL_1(P2_Set_ILDddlnnl_HL_1),
        .P2_Set_ILDddlnnl_SP_1(P2_Set_ILDddlnnl_SP_1),
        .P2_Set_ILDIXlnnl_0(P2_Set_ILDIXlnnl_0),
        .P2_Set_ILDIXlnnl_1(P2_Set_ILDIXlnnl_1),
        .P2_Set_ILDIYlnnl_0(P2_Set_ILDIYlnnl_0),
        .P2_Set_ILDIYlnnl_1(P2_Set_ILDIYlnnl_1),
        .P2_Set_ILDlnnlHL_0(P2_Set_ILDlnnlHL_0),
        .P2_Set_ILDlnnlHL_1(P2_Set_ILDlnnlHL_1),
        .P2_Set_ILDlnnldd_BC_0(P2_Set_ILDlnnldd_BC_0),
        .P2_Set_ILDlnnldd_DE_0(P2_Set_ILDlnnldd_DE_0),
        .P2_Set_ILDlnnldd_HL_0(P2_Set_ILDlnnldd_HL_0),
        .P2_Set_ILDlnnldd_SP_0(P2_Set_ILDlnnldd_SP_0),
        .P2_Set_ILDlnnldd_BC_1(P2_Set_ILDlnnldd_BC_1),
        .P2_Set_ILDlnnldd_DE_1(P2_Set_ILDlnnldd_DE_1),
        .P2_Set_ILDlnnldd_HL_1(P2_Set_ILDlnnldd_HL_1),
        .P2_Set_ILDlnnldd_SP_1(P2_Set_ILDlnnldd_SP_1),
        .P2_Set_ILDlnnlIX_0(P2_Set_ILDlnnlIX_0),
        .P2_Set_ILDlnnlIX_1(P2_Set_ILDlnnlIX_1),
        .P2_Set_ILDlnnlIY_0(P2_Set_ILDlnnlIY_0),
        .P2_Set_ILDlnnlIY_1(P2_Set_ILDlnnlIY_1),
        .P2_Set_IADDAn(P2_Set_IADDAn),
        .P2_Set_IADDAlIXtdl(P2_Set_IADDAlIXtdl),
        .P2_Set_IADDAlIYtdl(P2_Set_IADDAlIYtdl),
        .P2_Set_IADCAn(P2_Set_IADCAn),
        .P2_Set_IADCAlIXtdl(P2_Set_IADCAlIXtdl),
        .P2_Set_IADCAlIYtdl(P2_Set_IADCAlIYtdl),
        .P2_Set_ISUBAn(P2_Set_ISUBAn),
        .P2_Set_ISUBAlIXtdl(P2_Set_ISUBAlIXtdl),
        .P2_Set_ISUBAlIYtdl(P2_Set_ISUBAlIYtdl),
        .P2_Set_ISBCAn(P2_Set_ISBCAn),
        .P2_Set_ISBCAlIXtdl(P2_Set_ISBCAlIXtdl),
        .P2_Set_ISBCAlIYtdl(P2_Set_ISBCAlIYtdl),
        .P2_Set_IANDn(P2_Set_IANDn),
        .P2_Set_IANDlIXtdl(P2_Set_IANDlIXtdl),
        .P2_Set_IANDlIYtdl(P2_Set_IANDlIYtdl),
        .P2_Set_IORn(P2_Set_IORn),
        .P2_Set_IORlIXtdl(P2_Set_IORlIXtdl),
        .P2_Set_IORlIYtdl(P2_Set_IORlIYtdl),
        .P2_Set_IXORn(P2_Set_IXORn),
        .P2_Set_IXORlIXtdl(P2_Set_IXORlIXtdl),
        .P2_Set_IXORlIYtdl(P2_Set_IXORlIYtdl),
        .P2_Set_ICPn(P2_Set_ICPn),
        .P2_Set_ICPlIXtdl(P2_Set_ICPlIXtdl),
        .P2_Set_ICPlIYtdl(P2_Set_ICPlIYtdl),
        .P2_Set_IINClIXtdl(P2_Set_IINClIXtdl),
        .P2_Set_IINClIYtdl(P2_Set_IINClIYtdl),
        .P2_Set_IDEClIXtdl(P2_Set_IDEClIXtdl),
        .P2_Set_IDEClIYtdl(P2_Set_IDEClIYtdl),
        .P2_Set_IJPnn_0(P2_Set_IJPnn_0),
        .P2_Set_IJPnn_1(P2_Set_IJPnn_1),
        .P2_Set_IJPccnn_0_0(P2_Set_IJPccnn_0_0),
        .P2_Set_IJPccnn_1_0(P2_Set_IJPccnn_1_0),
        .P2_Set_IJPccnn_2_0(P2_Set_IJPccnn_2_0),
        .P2_Set_IJPccnn_3_0(P2_Set_IJPccnn_3_0),
        .P2_Set_IJPccnn_4_0(P2_Set_IJPccnn_4_0),
        .P2_Set_IJPccnn_5_0(P2_Set_IJPccnn_5_0),
        .P2_Set_IJPccnn_6_0(P2_Set_IJPccnn_6_0),
        .P2_Set_IJPccnn_7_0(P2_Set_IJPccnn_7_0),
        .P2_Set_IJPccnn_0_1(P2_Set_IJPccnn_0_1),
        .P2_Set_IJPccnn_1_1(P2_Set_IJPccnn_1_1),
        .P2_Set_IJPccnn_2_1(P2_Set_IJPccnn_2_1),
        .P2_Set_IJPccnn_3_1(P2_Set_IJPccnn_3_1),
        .P2_Set_IJPccnn_4_1(P2_Set_IJPccnn_4_1),
        .P2_Set_IJPccnn_5_1(P2_Set_IJPccnn_5_1),
        .P2_Set_IJPccnn_6_1(P2_Set_IJPccnn_6_1),
        .P2_Set_IJPccnn_7_1(P2_Set_IJPccnn_7_1),
        .P2_Set_IJRe(P2_Set_IJRe),
        .P2_Set_IJRCe(P2_Set_IJRCe),
        .P2_Set_IJRNCe(P2_Set_IJRNCe),
        .P2_Set_IJRZe(P2_Set_IJRZe),
        .P2_Set_IJRNZe(P2_Set_IJRNZe),
        .P2_Set_IDJNZe(P2_Set_IDJNZe),
        .P2_Set_ICALLnn_0(P2_Set_ICALLnn_0),
        .P2_Set_ICALLnn_1(P2_Set_ICALLnn_1),
        .P2_Set_ICALLnn_0_0(P2_Set_ICALLccnn_0_0),
        .P2_Set_ICALLnn_1_0(P2_Set_ICALLccnn_1_0),
        .P2_Set_ICALLnn_2_0(P2_Set_ICALLccnn_2_0),
        .P2_Set_ICALLnn_3_0(P2_Set_ICALLccnn_3_0),
        .P2_Set_ICALLnn_4_0(P2_Set_ICALLccnn_4_0),
        .P2_Set_ICALLnn_5_0(P2_Set_ICALLccnn_5_0),
        .P2_Set_ICALLnn_6_0(P2_Set_ICALLccnn_6_0),
        .P2_Set_ICALLnn_7_0(P2_Set_ICALLccnn_7_0),
        .P2_Set_ICALLnn_0_1(P2_Set_ICALLccnn_0_1),
        .P2_Set_ICALLnn_1_1(P2_Set_ICALLccnn_1_1),
        .P2_Set_ICALLnn_2_1(P2_Set_ICALLccnn_2_1),
        .P2_Set_ICALLnn_3_1(P2_Set_ICALLccnn_3_1),
        .P2_Set_ICALLnn_4_1(P2_Set_ICALLccnn_4_1),
        .P2_Set_ICALLnn_5_1(P2_Set_ICALLccnn_5_1),
        .P2_Set_ICALLnn_6_1(P2_Set_ICALLccnn_6_1),
        .P2_Set_ICALLnn_7_1(P2_Set_ICALLccnn_7_1),
        .P2_Set_IINAlnl(P2_Set_IINAlnl),
        .P2_Set_IOUTlnlA(P2_Set_IOUTlnlA),
        .P2_Reset_ITABLE(P2_Reset_ITABLE),
        .P2_Reset_ALLUNOFFICIALFF(P2_Reset_ALL_except_CRESET),
        .notIFF1(notIFF1),
        .IFF2(IFF2),
        .IMFa(IMFa),
        .IMFb(IMFb),
        .TINT(TINT),
        .TNMI(TNMI),
        .TRESET(TRESET),
        .TWAIT(TWAIT),
        .notLHALT(notLHALT),
        .notCM1(notCM1),
        .notCMR(notCMR),
        .notCMA(notCMA),
        .notCBUSRQ(notCBUSRQ),
        .notCRESET(notCRESET),
        .notCNMI(notCNMI),
        .notCINT0(notCINT0),
        .notCINT0_RST(notCINT0_RST),
        .notCINT0_CALL(notCINT0_CALL),
        .notCINT1(notCINT1),
        .notCINT2(notCINT2),
        .XIX(XIX),
        .XIX4_0(XIX4_0),
        .XIX4_1(XIX4_1),
        .XIY(XIY),
        .XIY4_0(XIY4_0),
        .XIY4_1(XIY4_1),
        .XOTR(XOTR),
        .XBIT(XBIT),
        .notXIX(notXIX),
        .notXIX4_0(notXIX4_0),
        .notXIX4_1(notXIX4_1),
        .notXIY(notXIY),
        .notXIY4_0(notXIY4_0),
        .notXIY4_1(notXIY4_1),
        .notXOTR(notXOTR),
        .notXBIT(notXBIT),
        .ITABLE(ITABLE),
        .notITABLE(notITABLE)
    );

    INTERFACE interface( // 952 + 37
        .notA(notA),
        .notF(notF),
        .notB(notB),
        .notC(notC),
        .notD(notD),
        .notE(notE),
        .notH(notH),
        .notL(notL),
        .notDt(notDt),
        .notDtex(notDtex),
        .notR(notR),
        .notI(notI),
        .notOP(notOP),
        .notOPold(notOPold),
        .notPC(notPC),
        .notSP(notSP),
        .notIX(notIX),
        .notIY(notIY),
        .notALU(notALU),
        // Ad
        .notPI_SelectAd_PC(~PI_SelectAd_PC),
        .notPI_SelectAd_SP(~PI_SelectAd_SP),
        .notPI_SelectAd_BC(~PI_SelectAd_BC),
        .notPI_SelectAd_DE(~PI_SelectAd_DE),
        .notPI_SelectAd_HL(~PI_SelectAd_HL),
        .notPI_SelectAd_IR(~PI_SelectAd_IR),
        .notPI_SelectAd_DtexDt(~PI_SelectAd_DtexDt),
        .notPI_SelectAd_OPOPold(~PI_SelectAd_OPOPold),
        .notPI_SelectAd_ALU(~PI_SelectAd_ALU),
        .notPI_SelectAd_AOP(~PI_SelectAd_AOP),
        .PI_SelectAdt1(PI_SelectAdt1),
        .notPI_Activate_Ad_high(~PI_Activate_Ad_high),
        .notPI_Activate_Ad_low(~PI_Activate_Ad_low),
        // Dt
        .notPI_SelectDt_PC_high(~PI_SelectDt_PC_high),
        .notPI_SelectDt_PC_low(~PI_SelectDt_PC_low),
        .notPI_SelectDt_IX_high(~PI_SelectDt_IX_high),
        .notPI_SelectDt_IX_low(~PI_SelectDt_IX_low),
        .notPI_SelectDt_IY_high(~PI_SelectDt_IY_high),
        .notPI_SelectDt_IY_low(~PI_SelectDt_IY_low),
        .notPI_SelectDt_A(~PI_SelectDt_A),
        .notPI_SelectDt_F(~PI_SelectDt_F),
        .notPI_SelectDt_B(~PI_SelectDt_B),
        .notPI_SelectDt_C(~PI_SelectDt_C),
        .notPI_SelectDt_D(~PI_SelectDt_D),
        .notPI_SelectDt_E(~PI_SelectDt_E),
        .notPI_SelectDt_H(~PI_SelectDt_H),
        .notPI_SelectDt_L(~PI_SelectDt_L),
        .notPI_SelectDt_OP(~PI_SelectDt_OP),
        .notPI_SelectDt_Dt(~PI_SelectDt_Dt),
        .notPI_SelectDt_Dtex(~PI_SelectDt_Dtex),
        .notPI_SelectDt_SP_low(~PI_SelectDt_SP_low),
        .notPI_SelectDt_SP_high(~PI_SelectDt_SP_high),
        .notPI_Activate_Dt(~PI_Activate_Dt),
        // out
        .notPI_Flag_BUSAK(~PI_Flag_BUSAK),
        .notPI_Flag_RFSH(~PI_Flag_RFSH),
        .notPI_Flag_M1(~PI_Flag_M1),
        .notPI_Flag_HALT(notLHALT),
        .PI_Nullify_MREQ(PI_Nullify_MREQ),
        .PI_Nullify_RD(PI_Nullify_RD),
        .PI_Nullify_WR(PI_Nullify_WR),
        .PI_Nullify_IORQ(PI_Nullify_IORQ),
        .notPI_Flag_MREQ(~PI_Flag_MREQ),
        .notPI_Flag_RD(~PI_Flag_RD),
        .notPI_Flag_WR(~PI_Flag_WR),
        .notPI_Flag_IORQ(~PI_Flag_IORQ),
        // interface
        .interfaceAd(interfaceAd),
        // 本当はinterfaceDt_inとinterfaceDt_outはinoutで同一だけどdigitalJSがエラーおこすので分けている
        .interfaceDt_in(interfaceDt_in),
        .interfaceDt_out(interfaceDt_out),
        .Din(Din),
        .interfaceBUSAK(interfaceBUSAK),
        .interfaceRFSH(interfaceRFSH),
        .interfaceM1(interfaceM1),
        .interfaceHALT(interfaceHALT),
        .interfaceMREQ(interfaceMREQ),
        .interfaceRD(interfaceRD),
        .interfaceWR(interfaceWR),
        .interfaceIORQ(interfaceIORQ)
    );

    REGISTER reg_( // 3834 + 34
        .Clk(Clk),
        .notClk(notClk),
        .notALUResult(notALU),
        .Din(Din),
        .notALULow0(notALULow0),
        .notALULow7(notALULow7),
        .notCY4(notCY4),
        .notCY8(notCY8),
        .CY12(CY12),
        .CY16(CY16),
        .notIs8bitEqual(notIs8bitEqual),
        .notIsResultLow0(notIsResultLow0),
        .isResult0(isResult0),
        .DAA_Flag_H(DAA_Flag_H),
        .IFF2(IFF2),
        .CINT(CINT),
        .is16bitEqual(is16bitEqual),
        .is8bitOverflow(is8bitOverflow),
        .notIs8bitEvenParity(notIs8bitEvenParity),
        .is16bitOverflow(is16bitOverflow),
        .PR_InvertIn(PR_InvertIn),
        // AF
        .PR_Write_A(PR_Write_A),
        .PR_Ex_AF_AF(PR_Ex_AF_AF),
        .PF_Write_S(PF_Write_S),
        .notPF_Select_S_bit7(~PF_Select_S_bit7),
        .notPF_Select_S_bit15(~PF_Select_S_bit15),
        .notPF_Select_S_bit23(~PF_Select_S_bit23),
        .PF_Write_Z(PF_Write_Z),
        .notPF_Select_Z_bit19(~PF_Select_Z_bit19),
        .notPF_Select_Z_bit21(~PF_Select_Z_bit21),
        .notPF_Select_Z_bit24(~PF_Select_Z_bit24),
        .notPF_Select_Z_bit34(~PF_Select_Z_bit34),
        .notPF_Select_Z_bit40(~PF_Select_Z_bit40),
        .notPF_Select_Z_bit41(~PF_Select_Z_bit41),
        .notPF_Select_Z_bit42(~PF_Select_Z_bit42),
        .notPF_Select_Z_bit43(~PF_Select_Z_bit43),
        .notPF_Select_Z_bit44(~PF_Select_Z_bit44),
        .notPF_Select_Z_bit45(~PF_Select_Z_bit45),
        .notPF_Select_Z_bit46(~PF_Select_Z_bit46),
        .notPF_Select_Z_bit47(~PF_Select_Z_bit47),
        .PF_Write_H(PF_Write_H),
        .PF_Select_H_bit17(PF_Select_H_bit17),
        .notPF_Select_H_bit21(~PF_Select_H_bit21),
        .notPF_Select_H_bit22(~PF_Select_H_bit22),
        .notPF_Select_H_bit28(~PF_Select_H_bit28),
        .notPF_Select_H_bit30(~PF_Select_H_bit30),
        .notPF_Select_H_bit31(~PF_Select_H_bit31),
        .notPF_Select_H_bit35(~PF_Select_H_bit35),
        .PF_Write_PV(PF_Write_PV),
        .notPF_Select_PV_bit18(~PF_Select_PV_bit18),
        .notPF_Select_PV_bit20(~PF_Select_PV_bit20),
        .notPF_Select_PV_bit25(~PF_Select_PV_bit25),
        .notPF_Select_PV_bit27(~PF_Select_PV_bit27),
        .notPF_Select_PV_bit33(~PF_Select_PV_bit33),
        .PF_Write_C(PF_Write_C),
        .PF_Select_C_bit17(PF_Select_C_bit17),
        .notPF_Select_C_bit23(~PF_Select_C_bit23),
        .notPF_Select_C_bit26(~PF_Select_C_bit26),
        .notPF_Select_C_bit29(~PF_Select_C_bit29),
        .notPF_Select_C_bit32(~PF_Select_C_bit32),
        .notPF_Select_C_bit36(~PF_Select_C_bit36),
        .notPF_Select_C_bit37(~PF_Select_C_bit37),
        .notPF_Select_C_bit38(~PF_Select_C_bit38),
        .PF_Select_C_bit0(PF_Select_C_bit0),
        .PF_Write_N(PF_Write_N),
        .PF_Select_N_bit17(PF_Select_N_bit17),
        .PR_Write_F(PR_Write_F),
        // BC
        .PR_Exx(PR_Exx),
        .PR_Write_B(PR_Write_B),
        .PR_Write_C(PR_Write_C),
        // DE
        .PR_EX_DE_HL(PR_EX_DE_HL),
        .PR_Write_D(PR_Write_D),
        .PR_Write_E(PR_Write_E),
        // HL
        .PR_Write_H(PR_Write_H),
        .PR_Write_L(PR_Write_L),
        // PC
        .PR_Write_PC_high(PR_Write_PC_high),
        .PR_Write_PC_low(PR_Write_PC_low),
        .PR_Inc_PC(PR_Inc_PC),
        // SP
        .PR_Write_SP_high(PR_Write_SP_high),
        .PR_Write_SP_low(PR_Write_SP_low),
        .PR_Inc_SP(PR_Inc_SP),
        .PR_Dec_SP(PR_Dec_SP),
        // IX
        .PR_Write_IX_high(PR_Write_IX_high),
        .PR_Write_IX_low(PR_Write_IX_low),
        // IY
        .PR_Write_IY_high(PR_Write_IY_high),
        .PR_Write_IY_low(PR_Write_IY_low),
        // I
        .PR_Write_I(PR_Write_I),
        // Dt
        .PR_Write_Dt(PR_Write_Dt),
        // Dtex
        .PR_Write_Dtex(PR_Write_Dtex),
        // Dtcs
        .PI_ReadDtcs(PI_ReadDtcs),
        // OP
        .PR_Write_OP(PR_Write_OP),
        // OPold
        .PR_SlideOP(PR_SlideOP),
        // R
        .PR_Write_R(PR_Write_R),
        .PR_Inc_R(PR_Inc_R),
        // XPT
        .PR_Reset_XPT(PR_Reset_XPT),
        .notPR_Halt_XPT(~PR_Halt_XPT),
        .notA(notA),
        .notF(notF),
        .notB(notB),
        .notC(notC),
        .notD(notD),
        .notE(notE),
        .notH(notH),
        .notL(notL),
        .notPC(notPC),
        .notSP(notSP),
        .notIX(notIX),
        .notIY(notIY),
        .notI(notI),
        .notDt(notDt),
        .notDtex(notDtex),
        .Dtcs(Dtcs),
        .notDtcs(notDtcs),
        .OP(OP),
        .notOP(notOP),
        .OPold(OPold),
        .notOPold(notOPold),
        .notR(notR),
        .XPT(XPT),
        .notXPT(notXPT)
    );

endmodule